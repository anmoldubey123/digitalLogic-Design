`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/11/2025 08:09:53 AM
// Design Name: 
// Module Name: tb_muxsm
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_muxsm;
reg clk;
reg reset;
reg [15:0] sw;
wire [3:0] an;
wire [6:0] sseg;


time_multiplexing_main u1(
.clk(clk), .reset(reset), .sw(sw), .an(an), .sseg(sseg)
    );
    
initial
begin    

clk = 0;
reset = 1;
sw [15:0] = 0000000000000000;

#40;

reset = 0;
sw [3:0] = 4'b0001;

#40;

sw [3:0] = 4'b0010;

#40;

sw [3:0] = 4'b0011;

#40;

sw [3:0] = 4'b0100;

#40;

sw [3:0] = 4'b0101;

#40;

sw [3:0] = 4'b0110;

#40;

sw[3:0] = 4'b0111;

#40;

sw[3:0] = 4'b1000;

#40;

sw[3:0] = 4'b1001;

#40;

sw[3:0] = 4'b1010;

#40;

sw[3:0] = 4'b1011;

#40;

sw[3:0] = 4'b1100;

#40;

sw[3:0] = 4'b1101;

#40;

sw[3:0] = 4'b1110;

#40;

sw[3:0] = 4'b1111;

#40;

sw[7:4] = 4'b0001;

#40;

sw[7:4] = 4'b0010;

#40;

sw[7:4] = 4'b0011;

#40;

sw[7:4] = 4'b0100;

#40;

sw[7:4] = 4'b0101;

#40;

sw[7:4] = 4'b0110;

#40;

sw[7:4] = 4'b0111;

#40;

sw[7:4] = 4'b1000;

#40;

sw[7:4] = 4'b1001;

#40;

sw[7:4] = 4'b1010;

#40;

sw[7:4] = 4'b1011;

#40;

sw[7:4] = 4'b1100;

#40;

sw[7:4] = 4'b1101;

#40;

sw[7:4] = 4'b1110;

#40;

sw[7:4] = 4'b1111;

#40

sw[11:8] = 4'b0001;

#40;

sw[11:8] = 4'b0010;

#40;

sw[11:8] = 4'b0011;

#40;

sw[11:8] = 4'b0100;

#40;

sw[11:8] = 4'b0101;

#40;

sw[11:8] = 4'b0110;

#40;

sw[11:8] = 4'b0111;

#40;

sw[11:8] = 4'b1000;

#40;

sw[11:8] = 4'b1001;

#40;

sw[11:8] = 4'b1010;

#40;

sw[11:8] = 4'b1011;

#40;

sw[11:8] = 4'b1100;

#40;

sw[11:8] = 4'b1101;

#40;

sw[11:8] = 4'b1110;

#40;

sw[11:8] = 4'b1111;

#40;

sw[15:12] = 4'b0001;

#40;

sw[15:12] = 4'b0010;

#40;

sw[15:12] = 4'b0011;

#40;

sw[15:12] = 4'b0100;

#40;

sw[15:12] = 4'b0101;

#40;

sw[15:12] = 4'b0110;

#40;

sw[15:12] = 4'b0111;

#40;

sw[15:12] = 4'b1000;

#40;

sw[15:12] = 4'b1001;

#40;

sw[15:12] = 4'b1010;

#40;

sw[15:12] = 4'b1011;

#40;

sw[15:12] = 4'b1100;

#0;

sw[15:12] = 4'b1101;

#40;

sw[15:12] = 4'b1110;

#40;

sw[15:12] = 4'b1111;

end 

always 
#5 clk = ~clk;

endmodule
